package vhdlGame {
  type SSD is array(6 downto 0) of std_logic;
  type SSDArray is array(natural range <>) of SSD;
}